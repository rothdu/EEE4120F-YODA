`include "./Constants/constants.v"

module Paralellizer (
    
);

endmodule