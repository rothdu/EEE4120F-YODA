// `include "./Constants/constants.v"
`include "./Paralellizer/paralellizer.v"
`include "./Encrypter/encrypter.v"
`include "./Collector/collector.vh"

module TestBench (
    
);

endmodule