`include "./Constants/constants.vh"

module Encrypter (
    
);

endmodule