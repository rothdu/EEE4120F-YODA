`define KEY_WIDTH 32 // width of the key
`define KEY_ROTATION_WIDTH 5 // width of the key rotation bus between Paralellizer and Encrypter
`define ENCRYPTER_WIDTH 32 // width of the bus between the Paralellizer and Encrypter, and the Encrypter and Collector. In multiples of 4.
`define NUM_ENCRYPTERS 4 // number of Encrypters