`include "./Constants/constants.v"

module Encrypter (
    
);

endmodule