module Paralellizer_tb (
    
);

endmodule