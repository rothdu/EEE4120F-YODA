`include "./Constants/constants.v"

module Collector (
    
);

endmodule