`include "./Constants/constants.vh"
`include "./Paralellizer/parallelizer.sv"
`include "./Encrypter/encrypter.sv"
`include "./Collector/collector.sv"

module TopLevel_tb (
    
);

endmodule